magic
tech sky130A
magscale 1 2
timestamp 1740675467
<< pwell >>
rect -201 -768 201 768
<< psubdiff >>
rect -165 698 -69 732
rect 69 698 165 732
rect -165 636 -131 698
rect 131 636 165 698
rect -165 -698 -131 -636
rect 131 -698 165 -636
rect -165 -732 -69 -698
rect 69 -732 165 -698
<< psubdiffcont >>
rect -69 698 69 732
rect -165 -636 -131 636
rect 131 -636 165 636
rect -69 -732 69 -698
<< xpolycontact >>
rect -35 170 35 602
rect -35 -602 35 -170
<< xpolyres >>
rect -35 -170 35 170
<< locali >>
rect -165 698 -69 732
rect 69 698 165 732
rect -165 636 -131 698
rect 131 636 165 698
rect -165 -698 -131 -636
rect 131 -698 165 -636
rect -165 -732 -69 -698
rect 69 -732 165 -698
<< viali >>
rect -19 187 19 584
rect -19 -584 19 -187
<< metal1 >>
rect -25 584 25 596
rect -25 187 -19 584
rect 19 187 25 584
rect -25 175 25 187
rect -25 -187 25 -175
rect -25 -584 -19 -187
rect 19 -584 25 -187
rect -25 -596 25 -584
<< properties >>
string FIXED_BBOX -148 -715 148 715
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.86 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 11.704k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
