magic
tech sky130A
magscale 1 2
timestamp 1740675467
<< pwell >>
rect -201 -1082 201 1082
<< psubdiff >>
rect -165 1012 -69 1046
rect 69 1012 165 1046
rect -165 950 -131 1012
rect 131 950 165 1012
rect -165 -1012 -131 -950
rect 131 -1012 165 -950
rect -165 -1046 -69 -1012
rect 69 -1046 165 -1012
<< psubdiffcont >>
rect -69 1012 69 1046
rect -165 -950 -131 950
rect 131 -950 165 950
rect -69 -1046 69 -1012
<< xpolycontact >>
rect -35 484 35 916
rect -35 -916 35 -484
<< xpolyres >>
rect -35 -484 35 484
<< locali >>
rect -165 1012 -69 1046
rect 69 1012 165 1046
rect -165 950 -131 1012
rect 131 950 165 1012
rect -165 -1012 -131 -950
rect 131 -1012 165 -950
rect -165 -1046 -69 -1012
rect 69 -1046 165 -1012
<< viali >>
rect -19 501 19 898
rect -19 -898 19 -501
<< metal1 >>
rect -25 898 25 910
rect -25 501 -19 898
rect 19 501 25 898
rect -25 489 25 501
rect -25 -501 25 -489
rect -25 -898 -19 -501
rect 19 -898 25 -501
rect -25 -910 25 -898
<< properties >>
string FIXED_BBOX -148 -1029 148 1029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 5.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 29.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
