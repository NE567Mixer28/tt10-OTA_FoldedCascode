** sch_path: /home/ttuser/FoldedCascode_OTA/xschem/untitled.sch
.subckt untitled IN+ IN- OUT VDD GND Vp Vp1 Vc1 Vc2 Vc3
*.PININFO IN+:I IN-:I OUT:O VDD:B GND:B Vp:B Vp1:B Vc1:B Vc2:B Vc3:B
XM1 D1 IN+ S S sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 m=5
XM2 D2 IN- S S sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 m=5
XM3 D1 Vc1 GND GND sky130_fd_pr__nfet_01v8 L=10 W=2 nf=1 m=1
XM4 D2 Vc1 GND GND sky130_fd_pr__nfet_01v8 L=10 W=2 nf=1 m=1
XM5 G Vc2 D1 GND sky130_fd_pr__nfet_01v8 L=2 W=3 nf=1 m=1
XM6 OUT Vc2 D2 GND sky130_fd_pr__nfet_01v8 L=2 W=3 nf=1 m=1
XM7 G Vc3 D9 D9 sky130_fd_pr__pfet_01v8 L=5 W=25 nf=1 m=1
XM8 OUT Vc3 D10 D10 sky130_fd_pr__pfet_01v8 L=5 W=25 nf=1 m=1
XM9 D9 G VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=30 nf=1 m=1
XM10 D10 G VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=30 nf=1 m=1
XM11 S Vp1 net1 VDD sky130_fd_pr__pfet_01v8 L=5 W=5 nf=1 m=1
XM12 net1 Vp VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=5 nf=1 m=1
.ends
.end
