magic
tech sky130A
magscale 1 2
timestamp 1740675467
<< nwell >>
rect -696 -719 696 719
<< pmos >>
rect -500 -500 500 500
<< pdiff >>
rect -558 488 -500 500
rect -558 -488 -546 488
rect -512 -488 -500 488
rect -558 -500 -500 -488
rect 500 488 558 500
rect 500 -488 512 488
rect 546 -488 558 488
rect 500 -500 558 -488
<< pdiffc >>
rect -546 -488 -512 488
rect 512 -488 546 488
<< nsubdiff >>
rect -660 649 -564 683
rect 564 649 660 683
rect -660 587 -626 649
rect 626 587 660 649
rect -660 -649 -626 -587
rect 626 -649 660 -587
rect -660 -683 -564 -649
rect 564 -683 660 -649
<< nsubdiffcont >>
rect -564 649 564 683
rect -660 -587 -626 587
rect 626 -587 660 587
rect -564 -683 564 -649
<< poly >>
rect -500 581 500 597
rect -500 547 -484 581
rect 484 547 500 581
rect -500 500 500 547
rect -500 -547 500 -500
rect -500 -581 -484 -547
rect 484 -581 500 -547
rect -500 -597 500 -581
<< polycont >>
rect -484 547 484 581
rect -484 -581 484 -547
<< locali >>
rect -660 649 -564 683
rect 564 649 660 683
rect -660 587 -626 649
rect 626 587 660 649
rect -500 547 -484 581
rect 484 547 500 581
rect -546 488 -512 504
rect -546 -504 -512 -488
rect 512 488 546 504
rect 512 -504 546 -488
rect -500 -581 -484 -547
rect 484 -581 500 -547
rect -660 -649 -626 -587
rect 626 -649 660 -587
rect -660 -683 -564 -649
rect 564 -683 660 -649
<< viali >>
rect -484 547 484 581
rect -546 -488 -512 488
rect 512 -488 546 488
rect -484 -581 484 -547
<< metal1 >>
rect -496 581 496 587
rect -496 547 -484 581
rect 484 547 496 581
rect -496 541 496 547
rect -552 488 -506 500
rect -552 -488 -546 488
rect -512 -488 -506 488
rect -552 -500 -506 -488
rect 506 488 552 500
rect 506 -488 512 488
rect 546 -488 552 488
rect 506 -500 552 -488
rect -496 -547 496 -541
rect -496 -581 -484 -547
rect 484 -581 496 -547
rect -496 -587 496 -581
<< properties >>
string FIXED_BBOX -643 -666 643 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
